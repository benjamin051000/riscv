module memory #(
    parameter int WIDTH = 32
) (
    input logic [WIDTH-1:0] addr, // TODO replace if not useful
    output logic [WIDTH-1:0] data
);

// TODO RAM and MMU

endmodule
